module interfaces

interface IdOwner {
	id int
}

struct User {
	id int
}
