module interface

interface IdOwner {
	id int
}

struct User {
	id int
}
