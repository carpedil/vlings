module movie_book

import readline { read_line }
import time

struct SeatBooking {}

fn (sb SeatBooking) check_bookings(seats [][]string) {
	println('正在为您查询该场次电影的预定状态...')
	println('从上到下为1~6排,从左至右为1~8座')

	println('============================================')
	for row in seats {
		println('  ${row}')
		time.sleep(100 * time.millisecond)
	}
	println('============================================')
}

fn (sb SeatBooking) book_seat(mut seats [][]string) ! {
	row := read_line('预订第几排的座位呢？请输入 1~6 之间的数字:\n')!
	colum := read_line('预订这一排的第几座呢？请输入 1~8 之间的数字:\n')!

	row_index := row.int() - 1
	colum_index := colum.int() - 1
	if seats[row_index][colum_index] == '○' {
		println('正在为您预订指定座位...')
		seats[colum_index][colum_index] = '●'
		println('预订成功！座位号：${row_index + 1}排${colum_index + 1}座')
	} else {
		println('这个座位已经被预订了哦')
	}
}

struct Movie {
	name   string
	symbol string
mut:
	seats [][]string
}

fn (m Movie) get_movies() []Movie {
	return [
		Movie{
			name: '泰坦尼克号'
			symbol: r'
			+==================== 泰坦尼克号 =====================+

		▄▄▄▄▄▪   ▄▄▄▄▄  ▄▄▄·   ▐ ▄ ▪      ▄▄· 
		•██   ██  •██   ▐█ ▀█  •█▌▐█  ██  ▐█ ▌▪
		▐█.▪ ▐█·  ▐█. ▪▄█▀▀█  ▐█▐▐▌  ▐█· ██ ▄▄
		▐█▌ ·▐█▌  ▐█▌· ▐█ ▪▐▌ ██▐█▌  ▐█▌ ▐███▌
		▀▀▀  ▀▀▀  ▀▀▀   ▀  ▀  ▀▀ █  ▪▀▀▀ ·▀▀▀ 

		+===================== Titanic =====================+'
			seats: [['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '●', '○', '○', '●'],
				['○', '○', '●', '○', '●', '○', '○', '○'],
				['○', '○', '●', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '○', '○', '●', '○'],
				['●', '○', '○', '○', '●', '●', '●', '●']]
		},
		Movie{
			name: '卡门'
			symbol: r'
			+======================= 卡门 =======================+

		▄█▄    ██   █▄▄▄▄ █▀▄▀█ ▄███▄      ▄   
		█▀ ▀▄  █ █  █  ▄▀ █ █ █ █▀   ▀      █  
		█   ▀  █▄▄█ █▀▀▌  █ ▄ █ ██▄▄    ██   █ 
		█▄  ▄▀ █  █ █  █  █   █ █▄   ▄▀ █ █  █ 
		▀███▀     █   █      █  ▀███▀   █  █ █ 
					█   ▀      ▀           █   ██ 
				▀                              

		+====================== Carmen =====================+'
			seats: [['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '●', '●', '○', '○', '●', '●'],
				['○', '○', '○', '○', '○', '○', '●', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '●', '○', '○', '○', '●']]
		},
		Movie{
			name: '机器人总动员'
			symbol: r'
			+==================== 机器人总动员 ===================+

		 ██   █▄▄▄▄ █▀▄▀█ ▄███▄      ▄   ▄█▄   
		 █ █  █  ▄▀ █ █ █ █▀   ▀      █  █▀ ▀▄ 
		 █▄▄█ █  ▌  █ ▄ █ ██▄▄    ██   █ █▄▄█▀ 
		 █  █ █  █  █   █ █▄   ▄▀ █ █  █ █▄  ▄▀
		    █   █      █  ▀█ ██ ▀   █  █ ▀███▀ █ 
					█   ▀      ▀           █   ██ 
				▀                              

		+====================== WALL·E =====================+'
			seats: [['●', '○', '○', '○', '○', '○', '○', '○'],
				['●', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '●', '○', '●', '○'],
				['○', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '○', '○', '●', '○', '○', '○'],
				['●', '●', '○', '○', '○', '●', '○', '○']]
		},
		Movie{
			name: '黑客帝国'
			symbol: r'
		+===================== 黑客帝国 =====================+

		________            __  ___      __       _     
		/_  __/ /_  ___     /  |/  /___ _/ /______(_)  __
		/ / / __ \\/ _ \\   / /|_/ / __ `/ __/ ___/ / |/_/
		/ / / / / /  __/  / /  / / /_/ / /_/ /  / />  <  
		/_/ /_/ /_/\\___/  /_/  /_/\\__,_/\\__/_/  /_/_/|_|  

		+==================== The Matrix ===================+'
			seats: [['○', '●', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '●', '●', '○', '○', '●'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '○', '○', '○', '○']]
		},
		Movie{
			name: '雨人'
			symbol: r'
		+====================== 雨人 =======================+

		,---      --   ,-  -   -             --    -   -  
		|  - \  / /\ \ |(||  \| | |\    /| / /\ \ |  \| | 
		/_  __/ /_  ___     /  |/  /___ _/ /______(_)  __
		|   (  |  __  || || ||  | (_)|/  ||  __  || ||  | 
		/_  __/ /_  ___     /  |/  /___ _/ /______(_)  __
		/_  __/ /_  ___     /  |/  /___ _/ /______(_)  __
			(__)         (__)     (__)   (__)        (__)     

		+===================== Rain Man ====================+'
			seats: [['○', '○', '○', '○', '●', '○', '○', '●'],
				['○', '○', '○', '●', '●', '○', '○', '○'],
				['○', '●', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '●', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○']]
		},
	]
}

fn test_check_bookings() ! {
	movie := Movie{}
	movie_list := movie.get_movies()
	println(movie_list.map(it.name))
	println('============================================')
	for index, val in movie_list {
		println('#${index + 1} -------------- ${val.name}')
	}
	println('============================================')
	mov_index := read_line('请输入您要预定的电影序号:')!

	valid_mov_idx := []int{len: movie_list.len, init: index}
	idx := mov_index.int() - 1

	println(idx in valid_mov_idx)

	mut movie_selected := movie.get_movies()[mov_index.int() - 1]

	// booking := SeatBooking{}

	// booking.check_bookings(movie_selected.seats)

	// booking.book_seat(mut movie_selected.seats)!
}
