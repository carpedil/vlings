module main

// import  vweb
// import json

// struct ApiData {
// 	vweb.Context 
// 	server_name string//服务名
// 	api_content string //	Api格式化后的内容。格式化后的内容可以是JSON或XML。应该在页面加载后立
// 	test_count int  // 测试次数，不太准确，但可以作为排序算法的参数。 有利于SNI
// }


// ['/api/save';post]
// pub fn (mut api ApiData) diff() vweb.Result {
// 	// body := json.decode(ApiData,api.req.data) or {
// 	// 	api.set_status(400,'')
// 	// 	return api.text('Failed to decode json, error: $err')
// 	//  }
// 	 // save data to db 

// 	return api.json('data saved ')
// }

