module movie_book

import readline { read_line }
import time

fn test_check_bookings() ! {
	movie := Movie{}
	movie_list := movie.get_movies()
	// println(movie_list.map(it.name))

	for {
		println('============================================')
		println('#场次\t\t电影名称')
		println('--------------------------------------------')

		for index, val in movie_list {
			println('#${index + 1} -------------- ${val.name}')
		}
		println('============================================')
		mov_index := read_line('请输入您要预定的电影场次: ')!

		valid_mov_idx := []int{len: movie_list.len, init: index}
		idx := mov_index.trim_space().int() - 1

		if idx >= 0 && idx < valid_mov_idx.len {
			mut movie_selected := movie.get_movies()[idx]
			println(movie_selected.symbol.trim_space())

			booking := SeatBooking{}

			booking.check_bookings(mut movie_selected.seats)!
		} else {
			println('请输入正确的电影场次: ')
		}
	}
}

struct SeatBooking {}

fn (sb SeatBooking) check_bookings(mut seats [][]string) ! {
	println('正在为您查询该场次电影的预定状态...')
	println('从上到下为1~6排,从左至右为1~8座')

	println('============================================')
	for row in seats {
		println('  ${row}')
		time.sleep(100 * time.millisecond)
	}
	println('============================================')
	sb.book_seat(mut seats)!
}

fn (sb SeatBooking) book_seat(mut seats [][]string) ! {
	row_label:
	row := read_line('预订第几排的座位呢？请输入 1~6 之间的数字: ')!

	row_index := row.trim_space().int() - 1
	if row_index >= 0 && row_index < 6 {
		colum_label:
		colum := read_line('预订这一排的第几座呢？请输入 1~8 之间的数字: ')!

		colum_index := colum.trim_space().int() - 1
		if colum_index >= 0 && colum_index < 8 {
			if seats[row_index][colum_index] == '○' {
				println('正在为您预订指定座位...')
				seats[row_index][colum_index] = '●'
				println('预订成功！座位号：${row_index + 1}排${colum_index + 1}座')
				time.sleep(3 * time.second)
				return
			} else {
				println('这个座位已经被预订了哦')
				return
			}
		} else {
			unsafe {
				println('输入有误! 请重新输入')
				goto colum_label
			}
		}
	} else {
		unsafe {
			println('输入有误! 请重新输入')
			goto row_label
		}
	}
}

struct Movie {
	name   string
	symbol string
mut:
	seats [][]string
}

fn (m Movie) get_movies() []Movie {
	return [
		Movie{
			name: '泰坦尼克号'
			symbol: r'
+==================== 泰坦尼克号 =====================+

  ▄▄▄▄▄▪   ▄▄▄▄▄  ▄▄▄·   ▐ ▄ ▪      ▄▄· 
  •██   ██  •██   ▐█ ▀█  •█▌▐█  ██  ▐█ ▌▪
  ▐█.▪ ▐█·  ▐█. ▪▄█▀▀█  ▐█▐▐▌  ▐█· ██ ▄▄
  ▐█▌ ·▐█▌  ▐█▌· ▐█ ▪▐▌ ██▐█▌  ▐█▌ ▐███▌
  ▀▀▀  ▀▀▀  ▀▀▀   ▀  ▀  ▀▀ █  ▪▀▀▀ ·▀▀▀ 

+===================== Titanic =====================+'
			seats: [['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '●', '○', '○', '●'],
				['○', '○', '●', '○', '●', '○', '○', '○'],
				['○', '○', '●', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '○', '○', '●', '○'],
				['●', '○', '○', '○', '●', '●', '●', '●']]
		},
		Movie{
			name: '卡门'
			symbol: r'
+======================= 卡门 =======================+

  ▄█▄    ██   █▄▄▄▄ █▀▄▀█ ▄███▄      ▄   
  █▀ ▀▄  █ █  █  ▄▀ █ █ █ █▀   ▀      █  
  █   ▀  █▄▄█ █▀▀▌  █ ▄ █ ██▄▄    ██   █ 
  █▄  ▄▀ █  █ █  █  █   █ █▄   ▄▀ █ █  █ 
  ▀███▀     █   █      █  ▀███▀   █  █ █ 
            █   ▀      ▀           █   ██ 
          ▀                              

+====================== Carmen =====================+'
			seats: [['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '●', '●', '○', '○', '●', '●'],
				['○', '○', '○', '○', '○', '○', '●', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '●', '○', '○', '○', '●']]
		},
		Movie{
			name: '机器人总动员'
			symbol: r"
+==================== 机器人总动员 ===================+

   (`\ .-') /`  ('-.                           ('-.   
    `.( OO ),' ( OO ).-.                     _(  OO)  
 ,--./  .--.   / . --. / ,--.      ,--.     (,------. 
 |      |  |   | \-.  \  |  |.-')  |  |.-')  |  .---' 
 |  |   |  |,.-'-'  |  | |  | OO ) |  | OO ) |  |     
 |  |.'.|  |_)\| |_.'  | |  |`-' | |  |`-' |(|  '--.  
 |         |   |  .-.  |(|  '---.'(|  '---.' |  .--'  
 |   ,'.   |   |  | |  | |      |  |      |  |  `---. 
 '--'   '--'   `--' `--' `------'  `------'  `------'  

+====================== WALL·E =====================+"
			seats: [['●', '○', '○', '○', '○', '○', '○', '○'],
				['●', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '●', '○', '●', '○'],
				['○', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '○', '○', '●', '○', '○', '○'],
				['●', '●', '○', '○', '○', '●', '○', '○']]
		},
		Movie{
			name: '黑客帝国'
			symbol: r'
+===================== 黑客帝国 =====================+

   ________            __  ___      __       _     
  /_  __/ /_  ___     /  |/  /___ _/ /______(_)  __
   / / / __ \/ _ \   / /|_/ / __ `/ __/ ___/ / |/_/
  / / / / / /  __/  / /  / / /_/ / /_/ /  / />  <  
 /_/ /_/ /_/\___/  /_/  /_/\__,_/\__/_/  /_/_/|_|  

+==================== The Matrix ===================+'
			seats: [['○', '●', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '●', '●', '○', '○', '●'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '●'],
				['○', '○', '●', '○', '○', '○', '○', '○']]
		},
		Movie{
			name: '雨人'
			symbol: r"
+====================== 雨人 =======================+

  ,---.    .--.  ,-..-. .-.           .--.  .-. .-. 
  | .-.\  / /\ \ |(||  \| | |\    /| / /\ \ |  \| | 
  | `-'/ / /__\ \(_)|   | | |(\  / |/ /__\ \|   | | 
  |   (  |  __  || || |\  | (_)\/  ||  __  || |\  | 
  | |\ \ | |  |)|| || | |)| | \  / || |  |)|| | |)| 
  |_| \)\|_|  (_)`-'/(  (_) | |\/| ||_|  (_)/(  (_) 
      (__)         (__)     '-'  '-'       (__)     

+===================== Rain Man ====================+"
			seats: [['○', '○', '○', '○', '●', '○', '○', '●'],
				['○', '○', '○', '●', '●', '○', '○', '○'],
				['○', '●', '○', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○'],
				['○', '○', '●', '○', '○', '○', '○', '○'],
				['○', '○', '○', '○', '○', '○', '○', '○']]
		},
	]
}
